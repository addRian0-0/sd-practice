library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Convertidores is 

	Port(
	
	);

end Convertidores;

architecture Ecuaciones of Convertidores is 

begin

end Ecuaciones;